library IEEE;
use IEEE.std_logic_1164.all;

entity clk_gen is
	port 
	(
		clk_in	:	in		std_logic;
		clk_out	:	out		std_logic
	);
end clk_gen;



architecture RTL of clk_gen is
begin


end RTL;